`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:03:08 11/22/2019 
// Design Name: 
// Module Name:    Pause_unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Pause_unit(
    input [31:0] IRD,
    input Clk,
    input Reset,
    output PauseD,
    output ClearE,
    output PauseF
    );


endmodule
